** sch_path: /home/gregu/gusharov_Analog_Bootcamp/analog/build/schematic/untitled.sch
**.subckt untitled
**.ends
.end
